
`timescale 1 ns / 1 ps
`timescale 1ns / 1ps
/*
```verilog
*/
// *******************************************************************************
// Company: Fpga Publish
// Engineer: FP 
// 
// Create Date: 2023/09/09 20:52:21
// Design Name: 
// Module Name: axi_cmd_v1_0
// Project Name: 
// Target Devices: ZYNQ7010 | XCZU2CG | Kintex7
// Tool Versions: 2021.1
// Description: 
//         * 
// Dependencies: 
//         * 
// Revision: 0.01 
// Revision 0.01 - File Created
//          1.1  - fix slaver not match error
// Additional Comments:
// 
// *******************************************************************************

	module axi_cmd_v1_0 #
	(
		// Users to add parameters here

		// User parameters ends
		// Do not modify the parameters beyond this line


		// Parameters of Axi Slave Bus Interface S00_AXI
		parameter integer C_S00_AXI_DATA_WIDTH	= 32,
		parameter integer C_S00_AXI_ADDR_WIDTH	= 9
	)
	(
		// Users to add ports here
        // Users to add ports here
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg0 ,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg1 ,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg2 ,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg3 ,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg4 ,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg5 ,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg6 ,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg7 ,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg8 ,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg9 ,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg10,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg11,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg12,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg13,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg14,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg15,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg16,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg17,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg18,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg19,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg20,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg21,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg22,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg23,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg24,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg25,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg26,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg27,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg28,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg29,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg30,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg31,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg32,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg33,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg34,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg35,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg36,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg37,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg38,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg39,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg40,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg41,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg42,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg43,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg44,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg45,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg46,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg47,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg48,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg49,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg50,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg51,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg52,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg53,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg54,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg55,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg56,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg57,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg58,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg59,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg60,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg61,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg62,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg63,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg64,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg65,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg66,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg67,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg68,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg69,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg70,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg71,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg72,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg73,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg74,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg75,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg76,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg77,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg78,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg79,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg80,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg81,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg82,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg83,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg84,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg85,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg86,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg87,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg88,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg89,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg90,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg91,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg92,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg93,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg94,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg95,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg96,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg97,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg98,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg99,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg100,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg101,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg102,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg103,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg104,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg105,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg106,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg107,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg108,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg109,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg110,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg111,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg112,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg113,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg114,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg115,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg116,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg117,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg118,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg119,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg120,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg121,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg122,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg123,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg124,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg125,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg126,
        output  [C_S00_AXI_DATA_WIDTH-1:0]    o_slv_reg127,
		// User ports ends
		// Do not modify the ports beyond this line


		// Ports of Axi Slave Bus Interface S00_AXI
		input wire  s00_axi_aclk,
		input wire  s00_axi_aresetn,
		input wire [C_S00_AXI_ADDR_WIDTH-1 : 0] s00_axi_awaddr,
		input wire [2 : 0] s00_axi_awprot,
		input wire  s00_axi_awvalid,
		output wire  s00_axi_awready,
		input wire [C_S00_AXI_DATA_WIDTH-1 : 0] s00_axi_wdata,
		input wire [(C_S00_AXI_DATA_WIDTH/8)-1 : 0] s00_axi_wstrb,
		input wire  s00_axi_wvalid,
		output wire  s00_axi_wready,
		output wire [1 : 0] s00_axi_bresp,
		output wire  s00_axi_bvalid,
		input wire  s00_axi_bready,
		input wire [C_S00_AXI_ADDR_WIDTH-1 : 0] s00_axi_araddr,
		input wire [2 : 0] s00_axi_arprot,
		input wire  s00_axi_arvalid,
		output wire  s00_axi_arready,
		output wire [C_S00_AXI_DATA_WIDTH-1 : 0] s00_axi_rdata,
		output wire [1 : 0] s00_axi_rresp,
		output wire  s00_axi_rvalid,
		input wire  s00_axi_rready
	);
// Instantiation of Axi Bus Interface S00_AXI
	axi_cmd_v1_0_S00_AXI # ( 
		.C_S_AXI_DATA_WIDTH(C_S00_AXI_DATA_WIDTH),
		.C_S_AXI_ADDR_WIDTH(C_S00_AXI_ADDR_WIDTH)
	) axi_cmd_v1_0_S00_AXI_inst (
        
        .o_slv_reg0     (o_slv_reg0  ),
        .o_slv_reg1     (o_slv_reg1  ),
        .o_slv_reg2     (o_slv_reg2  ),
        .o_slv_reg3     (o_slv_reg3  ),
        .o_slv_reg4     (o_slv_reg4  ),
        .o_slv_reg5     (o_slv_reg5  ),
        .o_slv_reg6     (o_slv_reg6  ),
        .o_slv_reg7     (o_slv_reg7  ),
        .o_slv_reg8     (o_slv_reg8  ),
        .o_slv_reg9     (o_slv_reg9  ),
        .o_slv_reg10    (o_slv_reg10 ),
        .o_slv_reg11    (o_slv_reg11 ),
        .o_slv_reg12    (o_slv_reg12 ),
        .o_slv_reg13    (o_slv_reg13 ),
        .o_slv_reg14    (o_slv_reg14 ),
        .o_slv_reg15    (o_slv_reg15 ),
        .o_slv_reg16    (o_slv_reg16 ),
        .o_slv_reg17    (o_slv_reg17 ),
        .o_slv_reg18    (o_slv_reg18 ),
        .o_slv_reg19    (o_slv_reg19 ),
        .o_slv_reg20    (o_slv_reg20 ),
        .o_slv_reg21    (o_slv_reg21 ),
        .o_slv_reg22    (o_slv_reg22 ),
        .o_slv_reg23    (o_slv_reg23 ),
        .o_slv_reg24    (o_slv_reg24 ),
        .o_slv_reg25    (o_slv_reg25 ),
        .o_slv_reg26    (o_slv_reg26 ),
        .o_slv_reg27    (o_slv_reg27 ),
        .o_slv_reg28    (o_slv_reg28 ),
        .o_slv_reg29    (o_slv_reg29 ),
        .o_slv_reg30    (o_slv_reg30 ),
        .o_slv_reg31    (o_slv_reg31 ),
        .o_slv_reg32    (o_slv_reg32 ),
        .o_slv_reg33    (o_slv_reg33 ),
        .o_slv_reg34    (o_slv_reg34 ),
        .o_slv_reg35    (o_slv_reg35 ),
        .o_slv_reg36    (o_slv_reg36 ),
        .o_slv_reg37    (o_slv_reg37 ),
        .o_slv_reg38    (o_slv_reg38 ),
        .o_slv_reg39    (o_slv_reg39 ),
        .o_slv_reg40    (o_slv_reg40 ),
        .o_slv_reg41    (o_slv_reg41 ),
        .o_slv_reg42    (o_slv_reg42 ),
        .o_slv_reg43    (o_slv_reg43 ),
        .o_slv_reg44    (o_slv_reg44 ),
        .o_slv_reg45    (o_slv_reg45 ),
        .o_slv_reg46    (o_slv_reg46 ),
        .o_slv_reg47    (o_slv_reg47 ),
        .o_slv_reg48    (o_slv_reg48 ),
        .o_slv_reg49    (o_slv_reg49 ),
        .o_slv_reg50    (o_slv_reg50 ),
        .o_slv_reg51    (o_slv_reg51 ),
        .o_slv_reg52    (o_slv_reg52 ),
        .o_slv_reg53    (o_slv_reg53 ),
        .o_slv_reg54    (o_slv_reg54 ),
        .o_slv_reg55    (o_slv_reg55 ),
        .o_slv_reg56    (o_slv_reg56 ),
        .o_slv_reg57    (o_slv_reg57 ),
        .o_slv_reg58    (o_slv_reg58 ),
        .o_slv_reg59    (o_slv_reg59 ),
        .o_slv_reg60    (o_slv_reg60 ),
        .o_slv_reg61    (o_slv_reg61 ),
        .o_slv_reg62    (o_slv_reg62 ),
        .o_slv_reg63    (o_slv_reg63 ),
        .o_slv_reg64    (o_slv_reg64 ),
        .o_slv_reg65    (o_slv_reg65 ),
        .o_slv_reg66    (o_slv_reg66 ),
        .o_slv_reg67    (o_slv_reg67 ),
        .o_slv_reg68    (o_slv_reg68 ),
        .o_slv_reg69    (o_slv_reg69 ),
        .o_slv_reg70    (o_slv_reg70 ),
        .o_slv_reg71    (o_slv_reg71 ),
        .o_slv_reg72    (o_slv_reg72 ),
        .o_slv_reg73    (o_slv_reg73 ),
        .o_slv_reg74    (o_slv_reg74 ),
        .o_slv_reg75    (o_slv_reg75 ),
        .o_slv_reg76    (o_slv_reg76 ),
        .o_slv_reg77    (o_slv_reg77 ),
        .o_slv_reg78    (o_slv_reg78 ),
        .o_slv_reg79    (o_slv_reg79 ),
        .o_slv_reg80    (o_slv_reg80 ),
        .o_slv_reg81    (o_slv_reg81 ),
        .o_slv_reg82    (o_slv_reg82 ),
        .o_slv_reg83    (o_slv_reg83 ),
        .o_slv_reg84    (o_slv_reg84 ),
        .o_slv_reg85    (o_slv_reg85 ),
        .o_slv_reg86    (o_slv_reg86 ),
        .o_slv_reg87    (o_slv_reg87 ),
        .o_slv_reg88    (o_slv_reg88 ),
        .o_slv_reg89    (o_slv_reg89 ),
        .o_slv_reg90    (o_slv_reg90 ),
        .o_slv_reg91    (o_slv_reg91 ),
        .o_slv_reg92    (o_slv_reg92 ),
        .o_slv_reg93    (o_slv_reg93 ),
        .o_slv_reg94    (o_slv_reg94 ),
        .o_slv_reg95    (o_slv_reg95 ),
        .o_slv_reg96    (o_slv_reg96 ),
        .o_slv_reg97    (o_slv_reg97 ),
        .o_slv_reg98    (o_slv_reg98 ),
        .o_slv_reg99    (o_slv_reg99 ),
        .o_slv_reg100   (o_slv_reg100),
        .o_slv_reg101   (o_slv_reg101),
        .o_slv_reg102   (o_slv_reg102),
        .o_slv_reg103   (o_slv_reg103),
        .o_slv_reg104   (o_slv_reg104),
        .o_slv_reg105   (o_slv_reg105),
        .o_slv_reg106   (o_slv_reg106),
        .o_slv_reg107   (o_slv_reg107),
        .o_slv_reg108   (o_slv_reg108),
        .o_slv_reg109   (o_slv_reg109),
        .o_slv_reg110   (o_slv_reg110),
        .o_slv_reg111   (o_slv_reg111),
        .o_slv_reg112   (o_slv_reg112),
        .o_slv_reg113   (o_slv_reg113),
        .o_slv_reg114   (o_slv_reg114),
        .o_slv_reg115   (o_slv_reg115),
        .o_slv_reg116   (o_slv_reg116),
        .o_slv_reg117   (o_slv_reg117),
        .o_slv_reg118   (o_slv_reg118),
        .o_slv_reg119   (o_slv_reg119),
        .o_slv_reg120   (o_slv_reg120),
        .o_slv_reg121   (o_slv_reg121),
        .o_slv_reg122   (o_slv_reg122),
        .o_slv_reg123   (o_slv_reg123),
        .o_slv_reg124   (o_slv_reg124),
        .o_slv_reg125   (o_slv_reg125),
        .o_slv_reg126   (o_slv_reg126),
        .o_slv_reg127   (o_slv_reg127),
        
		.S_AXI_ACLK(s00_axi_aclk),
		.S_AXI_ARESETN(s00_axi_aresetn),
		.S_AXI_AWADDR(s00_axi_awaddr),
		.S_AXI_AWPROT(s00_axi_awprot),
		.S_AXI_AWVALID(s00_axi_awvalid),
		.S_AXI_AWREADY(s00_axi_awready),
		.S_AXI_WDATA(s00_axi_wdata),
		.S_AXI_WSTRB(s00_axi_wstrb),
		.S_AXI_WVALID(s00_axi_wvalid),
		.S_AXI_WREADY(s00_axi_wready),
		.S_AXI_BRESP(s00_axi_bresp),
		.S_AXI_BVALID(s00_axi_bvalid),
		.S_AXI_BREADY(s00_axi_bready),
		.S_AXI_ARADDR(s00_axi_araddr),
		.S_AXI_ARPROT(s00_axi_arprot),
		.S_AXI_ARVALID(s00_axi_arvalid),
		.S_AXI_ARREADY(s00_axi_arready),
		.S_AXI_RDATA(s00_axi_rdata),
		.S_AXI_RRESP(s00_axi_rresp),
		.S_AXI_RVALID(s00_axi_rvalid),
		.S_AXI_RREADY(s00_axi_rready)
	);

	// Add user logic here

	// User logic ends

	endmodule
